// fc2__packed_params__packed_params_bias
localparam signed [7:0] fc2__packed_params__packed_params_bias [0:1] = '{
8'd0, 8'd0
};
