// fc1_zero_point
localparam signed [7:0] fc1_zero_point [0:0] = '{
8'd0
};
