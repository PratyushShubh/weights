// fc1_scale
localparam signed [7:0] fc1_scale [0:0] = '{
8'd1
};
