// fc2_zero_point
localparam signed [7:0] fc2_zero_point [0:0] = '{
8'd0
};
