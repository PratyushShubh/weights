// fc2_scale
localparam signed [7:0] fc2_scale [0:0] = '{
8'd1
};
